module game(input rst,clk, sel,next,output [1:0] a,b,c,d,e,f,g,h,i);


	


endmodule 